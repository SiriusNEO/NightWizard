module LS_EX (

);



endmodule