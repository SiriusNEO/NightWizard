module LSQueue (

);

endmodule