module LS_Executor (

);



endmodule