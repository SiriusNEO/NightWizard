module Fetcher(

);



endmodule