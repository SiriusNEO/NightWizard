// RISCV32I CPU top module
// port modification allowed for debugging purposes

`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/defines.v"

`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/if_unit/Fetcher.v"
`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/if_unit/PcReg.v"

`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/id_unit/Dispatcher.v"
`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/id_unit/Decoder.v"

`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/ex_unit/RS.v"
`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/ex_unit/RS_EX.v"

`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/pub_unit/MemCtrl.v"
`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/pub_unit/RegFile.v"
`include "/mnt/c/Users/17138/Desktop/CPU/NightWizard/cpu/src/pub_unit/ReOrderBuffer.v"

module cpu(
  input  wire                 clk_in,			// system clock signal
  input  wire                 rst_in,			// reset signal
	input  wire					        rdy_in,			// ready signal, pause cpu when low

  input  wire [ 7:0]          mem_din,		// data input bus
  output wire [ 7:0]          mem_dout,		// data output bus
  output wire [31:0]          mem_a,			// address bus (only 17:0 is used)
  output wire                 mem_wr,			// write/read signal (1 for write)
	
	input  wire                 io_buffer_full, // 1 if uart buffer is full
	
	output wire [31:0]			dbgreg_dout		// cpu register output (debugging demo)
);

// implementation goes here

// Specifications:
// - Pause cpu(freeze pc, registers, etc.) when rdy_in is low
// - Memory read result will be returned in the next cycle. Write takes 1 cycle(no need to wait)
// - Memory is of size 128KB, with valid address ranging from 0x0 to 0x20000
// - I/O port is mapped to address higher than 0x30000 (mem_a[17:16]==2'b11)
// - 0x30000 read: read a byte from input
// - 0x30000 write: write a byte to output (write 0x00 is ignored)
// - 0x30004 read: read clocks passed since cpu starts (in dword, 4 bytes)
// - 0x30004 write: indicates program stop (will output '\0' through uart tx)

// fetcher and memctrl
wire [`ADDR_LEN - 1 : 0] pc_if_mc;
wire [`INS_LEN - 1 : 0] inst_mc_if;
wire ena_if_mc, ok_flag_mc_if;

// fetcher and dispatcher
wire [`INS_LEN - 1 : 0] inst_if_dsp;
wire [`ADDR_LEN - 1 : 0] pc_if_dsp;
wire ok_flag_if_dsp;

// fetcher and pcreg
wire upd_if_pcr;
wire [`ADDR_LEN - 1 : 0] pc_pcr_if;

// full signal to fetcher
wire full_rs_if, full_lsb_if, full_rob_if;

// fetcher and decoder
wire [`INS_LEN - 1 : 0] inst_if_dcd;

// dispatcher and decoder
wire [`OPENUM_LEN - 1 : 0] openum_dcd_dsp;
wire [`REG_LEN - 1 : 0] rd_dcd_dsp, rs1_dcd_dsp, rs2_dcd_dsp;
wire [`DATA_LEN - 1 : 0] imm_dcd_dsp;

// dispatcher and rs
wire ena_dsp_rs;
wire [`OPENUM_LEN - 1 : 0] openum_dsp_rs;
wire [`DATA_LEN -1 : 0] V1_dsp_rs;
wire [`DATA_LEN -1 : 0] V2_dsp_rs;
wire [`ROB_LEN : 0] Q1_dsp_rs;
wire [`ROB_LEN : 0] Q2_dsp_rs;
wire [`ADDR_LEN -1 : 0] pc_dsp_rs;
wire [`ADDR_LEN -1 : 0] imm_dsp_rs;
wire [`ROB_LEN : 0] rob_id_dsp_rs;

// dispatcher and lsbuffer
wire ena_dsp_lsb;
wire [`OPENUM_LEN - 1 : 0] openum_dsp_lsb;
wire [`DATA_LEN -1 : 0] V1_dsp_lsb;
wire [`DATA_LEN -1 : 0] V2_dsp_lsb;
wire [`ROB_LEN : 0] Q1_dsp_lsb;
wire [`ROB_LEN : 0] Q2_dsp_lsb;
wire [`ADDR_LEN -1 : 0] imm_dsp_lsb;
wire [`ROB_LEN : 0] rob_id_dsp_lsb;

// dispatcher and rob
wire ena_dsp_rob;
wire [`REG_LEN - 1 : 0] rd_dsp_rob;
wire [`DATA_LEN - 1 : 0] data_dsp_rob;
wire [`ADDR_LEN - 1 : 0] pc_dsp_rob;
wire [`ROB_LEN : 0] rob_id_rob_dsp;

// dispatcher and regfile
wire [`REG_LEN - 1 : 0] rs1_dsp_reg;
wire [`REG_LEN - 1 : 0] rs2_dsp_reg;
wire [`DATA_LEN -1 : 0] V1_reg_dsp;
wire [`DATA_LEN -1 : 0] V2_reg_dsp;
wire [`ROB_LEN : 0] Q1_reg_dsp;
wire [`ROB_LEN : 0] Q2_reg_dsp;

// regfile and rob
wire [`ROB_LEN : 0] Q1_reg_rob;
wire [`ROB_LEN : 0] Q2_reg_rob;
wire Q1_ready_rob_reg;
wire Q2_ready_rob_reg;

// commit
// rob to reg
wire [`REG_LEN - 1 : 0] rd_rob_reg;
wire [`ROB_LEN : 0] Q_rob_reg;
wire [`DATA_LEN - 1 : 0] V_rob_reg;

// rs and rs_ex
wire [`OPENUM_LEN - 1 : 0] openum_rs_ex;
wire [`DATA_LEN - 1 : 0] V1_rs_ex;
wire [`DATA_LEN - 1 : 0] V2_rs_ex;
wire [`DATA_LEN - 1 : 0] imm_rs_ex;
wire [`ADDR_LEN - 1 : 0] pc_rs_ex;

// ls and ls_ex

// cdb
wire [`ROB_LEN : 0] rob_id_cdb;
wire [`DATA_LEN - 1 : 0] result_cdb;
wire [`ADDR_LEN - 1 : 0] target_pc_cdb;

PcReg pcReg(
  .rst(rst_in),
  .update(upd_if_pcr),
  .pc(pc_pcr_if)
);

Fetcher fetcher(
  .clk(clk_in),
  .rst(rst_in),
  .rdy(rdy_in),

  .inst_to_dcd(inst_if_dcd),

  .pc_to_mc(pc_if_mc),
  .ena_to_mc(ena_if_mc),

  .ok_flag_from_mc(ok_flag_mc_if),
  .inst_from_mc(inst_mc_if),

  .inst_to_dsp(inst_if_dsp),
  .pc_to_dsp(pc_if_dsp),
  .ok_flag_to_dsp(ok_flag_if_dsp),

  .pc_from_pcr(pc_pcr_if),
  .upd_to_pcr(upd_if_pcr)
);

Dispatcher dispatcher(
  .clk(clk_in),
  .rst(rst_in),
  .rdy(rdy_in),

  .ok_flag_from_if(ok_flag_if_dsp),
  .inst_from_if(inst_if_dsp),
  .pc_from_if(pc_if_dsp),

  // decoder
  .openum_from_dcd(openum_dcd_dsp),
  .rd_from_dcd(rd_dcd_dsp),
  .rs1_from_dcd(rs1_dcd_dsp),
  .rs2_from_dcd(rs2_dcd_dsp),
  .imm_from_dcd(imm_dcd_dsp),

  // to rob
  .ena_to_rob(ena_dsp_rob),
  .rd_to_rob(rd_dsp_rob),
  .pc_to_rob(pc_dsp_rob),
  // from rob
  .rob_id_from_rob(rob_id_rob_dsp),

  // to reg
  .rs1_to_reg(rs1_dsp_reg),
  .rs2_to_reg(rs2_dsp_reg), 
  // from reg
  .V1_from_reg(V1_reg_dsp),
  .V2_from_reg(V2_reg_dsp),
  .Q1_from_reg(Q1_reg_dsp),
  .Q2_from_reg(Q2_reg_dsp),

  // to rs
  .ena_to_rs(ena_dsp_rs),
  .openum_to_rs(openum_dsp_rs),
  .V1_to_rs(V1_dsp_rs),
  .V2_to_rs(V2_dsp_rs),
  .Q1_to_rs(Q1_dsp_rs),
  .Q2_to_rs(Q2_dsp_rs),
  .pc_to_rs(pc_dsp_rs),
  .imm_to_rs(imm_dsp_rs),
  .rob_id_to_rs(rob_id_dsp_rs),

  // to ls
  .openum_to_lsb(openum_dsp_lsb),
  .V1_to_lsb(V1_dsp_lsb),
  .V2_to_lsb(V2_dsp_lsb),
  .Q1_to_lsb(Q1_dsp_lsb),
  .Q2_to_lsb(Q2_dsp_lsb),
  .imm_to_lsb(imm_dsp_lsb),
  .rob_id_to_lsb(rob_id_dsp_lsb)
);

Decoder decoder(
  .ena(rdy_in),

  .inst(inst_if_dcd),

  .openum(openum_dcd_dsp),
  .rd(rd_dcd_dsp),
  .rs1(rs1_dcd_dsp),
  .rs2(rs2_dcd_dsp),
  .imm(imm_dcd_dsp)
);

RS rs(
  .clk(clk_in),
  .rst(rst_in),

  // from dsp
  .ena_from_dsp(ena_dsp_rs),
  .openum_from_dsp(openum_dsp_rs),
  .V1_from_dsp(V1_dsp_rs),
  .V2_from_dsp(V2_dsp_rs),
  .Q1_from_dsp(Q1_dsp_rs),
  .Q2_from_dsp(Q2_dsp_rs),
  .pc_from_dsp(pc_dsp_rs),
  .imm_from_dsp(imm_dsp_rs),
  .rob_id_from_dsp(rob_id_dsp_rs),

  // to ex
  .openum_to_ex(openum_rs_ex),
  .V1_to_ex(V1_rs_ex),
  .V2_to_ex(V2_rs_ex),
  .pc_to_ex(pc_rs_ex),
  .imm_to_ex(imm_rs_ex),

  // to cdb
  .rob_id_to_cdb(rob_id_cdb)
);

RS_EX rs_ex(
  .openum(openum_rs_ex),
  .V1(V1_rs_ex),
  .V2(V2_rs_ex),
  .imm(imm_rs_ex),
  .pc(pc_rs_ex),
  
  .result(result_cdb),
  .target_pc(target_pc_cdb)
);

ReOrderBuffer reOrderBuffer(
  .clk(clk_in),
  .rst(rst_in),

  // reply to reg_ready query
  // from reg
  .Q1_from_reg(Q1_reg_rob),
  .Q2_from_reg(Q2_reg_rob),
  // to reg
  .Q1_ready_to_reg(Q1_ready_rob_reg),
  .Q2_ready_to_reg(Q2_ready_rob_reg),

  // dsp allocate to rob
  // from dsp
  .ena_from_dsp(ena_dsp_rob),
  .rd_from_dsp(rd_dsp_rob),
  .pc_from_dsp(pc_dsp_rob),
  // to dsp
  .rob_id_to_dsp(rob_id_rob_dsp),

  // update rob by cdb
  // from cdb
  .rob_id_from_cdb(rob_id_cdb),
  .result_from_cdb(result_cdb),

  // commit
  // to reg
  .rd_to_reg(rd_rob_reg),
  .Q_to_reg(Q_rob_reg),
  .V_to_reg(V_rob_reg)
);

MemCtrl memCtrl(
  .clk(clk_in),
  .rst(rst_in),
  .rdy(rdy_in),

  // with ram
  .uart_full_from_ram(io_buffer_full),
  .wr_flag_to_ram(mem_wr),

  .addr_to_ram(mem_a),
    
  .data_i_from_ram(mem_din),
  .data_o_to_ram(mem_dout),

  // with fetcher
  .pc_from_if(pc_if_mc),
  .ena_from_if(ena_if_mc),
  .ok_flag_to_if(ok_flag_mc_if),
  .inst_to_if(inst_mc_if)
);

RegFile regFile(
  .clk(clk_in),
  .rst(rst_in),

  // from dsp
  .rs1_from_dsp(rs1_dsp_reg),
  .rs2_from_dsp(rs2_dsp_reg),

  // to dsp
  .V1_to_dsp(V1_reg_dsp),
  .V2_to_dsp(V2_reg_dsp),
  .Q1_to_dsp(Q1_reg_dsp),
  .Q2_to_dsp(Q2_reg_dsp),

  // to rob
  .Q1_to_rob(Q1_reg_rob),
  .Q2_to_rob(Q2_reg_rob),
  
  // from rob
  .Q1_ready_from_rob(Q1_ready_rob_reg),
  .Q2_ready_from_rob(Q2_ready_rob_reg)
);

always @(posedge clk_in)
  begin
    if (rst_in)
      begin
      
      end
    else if (!rdy_in)
      begin
      
      end
    else
      begin
      
      end
  end

endmodule